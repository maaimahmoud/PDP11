LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

package mine is
	
	type genericArrayofVector16bit is array (natural range <>) of std_logic_vector(15 downto 0);

	-- type genericArray is array (natural range <>) of std_logic_vector (15 downto 0);

end mine;


-- Package Body Section
package body mine is

	
end mine;


